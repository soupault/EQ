module filter (
	input wire [] 
	
	input wire i_rst_n,
	input wire i_clk,
	input wire i_ena,

	output reg [x:x] ,
	output reg x
);

always @(posedge i_clk or negedge i_rst_n)
begin
	if (~i_rst_n) begin
		
	end else begin
		
	end
end

endmodule
