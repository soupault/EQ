interface dut_if();

  logic clk;
  logic nrst;
  logic spdif;

endinterface: dut_if

