package my_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
// configuration object between TB and UVM
`include "my_dut_config.svh"
`include "my_transaction.svh"
`include "my_sequence.svh"
`include "my_sequencer.svh"
`include "my_driver.svh"
`include "my_monitor.svh"
`include "my_subscriber.svh"
`include "my_agent.svh"
`include "my_env.svh"
`include "my_test.svh"

endpackage: my_pkg

