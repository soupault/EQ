
`define AUX_SAMPLE    3:0
`define AUDIO_SAMPLE  23:4
`define VALIDITY      24
`define USER_DATA     25
`define CHNL_STATUS   26
`define PARITY        27

